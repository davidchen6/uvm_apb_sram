`ifndef APB_GLOBAL_PKG__SV
`define APB_GLOBAL_PKG__SV

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File Name: apb_global_pkg.sv
// Author: CCW
// Email: chengjiuweiye8@163.com
// Revision: 0.1
// Description: global package for holding global defines
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

package apb_global_pkg;
	//include global defines
	`include "tbf_defines.sv"

endpackage
`endif

